module top_gen_overlapped (clk, res_n, D1, D2, D3, F0, F1);
									
input logic 		 clk, res_n;
input logic [15:0] D1, D2, D3;
output logic			  F0, F1;

gen_overlapped UUT (clk, res_n, D1, D2, D3, F0, F1);

endmodule
