module debouncer (clk, inp, _rst)

input logic ;
output logic ;