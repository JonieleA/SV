module num2 (clk, rb, comb, out);

input logic clk, rb;
input logic [5:0] comb;
output logic out;
logic [48:0] w;
//Подключим делители
div #(.C(384_615)) DUT1(.clk(clk), .rb(rb), .out(w[0]));//65.41 Гц С большая октава
div #(.C(192_307)) DUT2(.clk(clk), .rb(rb), .out(w[1]));//130Гц С малая октава
div #(.C(95_419)) DUT3(.clk(clk), .rb(rb), .out(w[2]));//262 Гц С первая октава
div #(.C(47_801)) DUT4(.clk(clk), .rb(rb), .out(w[3]));//523 Гц С вторая октава
div #(.C(23_877)) DUT5(.clk(clk), .rb(rb), .out(w[4]));//1047 Гц С третья октава
div #(.C(11_944)) DUT6(.clk(clk), .rb(rb), .out(w[5]));//2093 Гц С четвёртая октава
div #(.C(5_958)) DUT7(.clk(clk), .rb(rb), .out(w[6]));//4196 Гц С пятая октава
div #(.C(337_837)) DUT8(.clk(clk), .rb(rb), .out(w[7]));//74 Гц D большая октава
div #(.C(168_918)) DUT9(.clk(clk), .rb(rb), .out(w[8]));//148 Гц D малая октава
div #(.C(85_034)) DUT10(.clk(clk), .rb(rb), .out(w[9]));//294 Гц D первая октава
div #(.C(42_589)) DUT11(.clk(clk), .rb(rb), .out(w[10]));//587 Гц D вторая октава
div #(.C(21_276)) DUT12(.clk(clk), .rb(rb), .out(w[11]));//1175 Гц D третья октава
div #(.C(10_642)) DUT13(.clk(clk), .rb(rb), .out(w[12]));//2349 Гц D четвёртая октава 
div #(.C(5_322)) DUT14(.clk(clk), .rb(rb), .out(w[13]));//4697 Гц D пятая октава
div #(.C(304_878)) DUT15(.clk(clk), .rb(rb), .out(w[14]));//82 Гц E большая октава
div #(.C(152_439)) DUT16(.clk(clk), .rb(rb), .out(w[15]));//164 Гц E малая октава
div #(.C(76_219)) DUT17(.clk(clk), .rb(rb), .out(w[16]));//328 Гц E первая октава
div #(.C(38_109)) DUT18(.clk(clk), .rb(rb), .out(w[17]));//656 Гц E вторая октава
div #(.C(19_054)) DUT19(.clk(clk), .rb(rb), .out(w[18]));//1312 Гц E третья октава
div #(.C(9_480)) DUT20(.clk(clk), .rb(rb), .out(w[19]));//2637 Гц E четвёртая октава
div #(.C(4_740)) DUT21(.clk(clk), .rb(rb), .out(w[20]));//5274 Гц E пятая октава
div #(.C(287_356)) DUT22(.clk(clk), .rb(rb), .out(w[21]));//87 Гц F большая октава
div #(.C(143_678)) DUT23(.clk(clk), .rb(rb), .out(w[22]));//174 Гц F малая октава
div #(.C(71_633)) DUT24(.clk(clk), .rb(rb), .out(w[23]));//349 Гц F первая октава
div #(.C(35_816)) DUT25(.clk(clk), .rb(rb), .out(w[24]));//698 Гц F вторая октава
div #(.C(17_908)) DUT26(.clk(clk), .rb(rb), .out(w[25]));//1396 Гц F третья октава
div #(.C(8_950)) DUT27(.clk(clk), .rb(rb), .out(w[26]));//2793 Гц F четвёртая октава
div #(.C(4_475)) DUT28(.clk(clk), .rb(rb), .out(w[27]));//5586 Гц F пятая октава
div #(.C(255_102)) DUT29(.clk(clk), .rb(rb), .out(w[28]));//98 Гц G большая октава
div #(.C(127_551)) DUT30(.clk(clk), .rb(rb), .out(w[29]));//196 Гц G малая октава
div #(.C(63_775)) DUT31(.clk(clk), .rb(rb), .out(w[30]));//392 Гц G первая октава
div #(.C(31_887)) DUT32(.clk(clk), .rb(rb), .out(w[31]));//784 Гц G вторая октава
div #(.C(15_943)) DUT33(.clk(clk), .rb(rb), .out(w[32]));//1568 Гц G третья октава
div #(.C(7_971)) DUT34(.clk(clk), .rb(rb), .out(w[33]));//3136 Гц G четвёртая октава
div #(.C(3_985)) DUT35(.clk(clk), .rb(rb), .out(w[34]));//6272 ГЦ G пятая октава
div #(.C(227_272)) DUT36(.clk(clk), .rb(rb), .out(w[35]));//110 Гц A большая октава
div #(.C(113_636)) DUT37(.clk(clk), .rb(rb), .out(w[36]));//220 Гц A малая октава
div #(.C(56_818)) DUT38(.clk(clk), .rb(rb), .out(w[37]));//440 Гц A первая октава
div #(.C(28_409)) DUT39(.clk(clk), .rb(rb), .out(w[38]));//880 Гц А вторая октава
div #(.C(14_204)) DUT40(.clk(clk), .rb(rb), .out(w[39]));//1760 Гц А третья октава
div #(.C(7_102)) DUT41(.clk(clk), .rb(rb), .out(w[40]));//3520 Гц А четвёртая октава
div #(.C(3_551)) DUT42(.clk(clk), .rb(rb), .out(w[41]));//7040 Гц А пятая октава
div #(.C(203_252)) DUT43(.clk(clk), .rb(rb), .out(w[42]));//123 Гц В большая октава
div #(.C(101_626)) DUT44(.clk(clk), .rb(rb), .out(w[43]));//246 Гц В малая октава
div #(.C(50_813)) DUT45(.clk(clk), .rb(rb), .out(w[44]));//492 Гц В первая октава
div #(.C(25_406)) DUT46(.clk(clk), .rb(rb), .out(w[45]));//984 Гц В вторая октава
div #(.C(12_703)) DUT47(.clk(clk), .rb(rb), .out(w[46]));//1968 Гц В третья октава
div #(.C(6_327)) DUT48(.clk(clk), .rb(rb), .out(w[47]));//3951 Гц В четвёртая октава
div #(.C(3_163)) DUT49(.clk(clk), .rb(rb), .out(w[48]));//7902 Гц В пятая октава

//От комбинации на выход передаётся сигнал соответствующего делителя				
always_comb begin
	case(comb)
	6'b000001 : out <= w[0] ;
	6'b001001 : out <= w[1] ;
	6'b010001 : out <= w[2] ;
	6'b011001 : out <= w[3] ;
	6'b100001 : out <= w[4] ;
	6'b101001 : out <= w[5] ;
	6'b110001 : out <= w[6] ;
	6'b000010 : out <= w[7] ;
	6'b001010 : out <= w[8] ;
	6'b010010 : out <= w[9] ;
	6'b011010 : out <= w[10] ;
	6'b100010 : out <= w[11] ;
	6'b101010 : out <= w[12] ;
   6'b110010 : out <= w[13] ;
	6'b000011 : out <= w[14] ;
	6'b001011 : out <= w[15] ;
	6'b010011 : out <= w[16] ;
	6'b011011 : out <= w[17] ;
	6'b100011 : out <= w[18] ;
	6'b101011 : out <= w[19] ;
	6'b110011 : out <= w[20] ;
	6'b000100 : out <= w[21] ;
	6'b001100 : out <= w[22] ;
	6'b010100 : out <= w[23] ;
	6'b011100 : out <= w[24] ;
	6'b100100 : out <= w[25] ;
	6'b101100 : out <= w[26] ;
	6'b110100 : out <= w[27] ;
	6'b000101 : out <= w[28] ;
	6'b001101 : out <= w[29] ;
	6'b010101 : out <= w[30] ;
	6'b011101 : out <= w[31] ;
	6'b100101 : out <= w[32] ;
   6'b101101 : out <= w[33] ;
	6'b110101 : out <= w[34] ;
	6'b000110 : out <= w[35] ;
	6'b001110 : out <= w[36] ;
	6'b010110 : out <= w[37] ;
	6'b011110 : out <= w[38] ;
	6'b100110 : out <= w[39] ;
	6'b101110 : out <= w[40] ;
	6'b110110 : out <= w[41] ;
	6'b000111 : out <= w[42] ;
   6'b001111 : out <= w[43] ;
	6'b010111 : out <= w[44] ;
	6'b011111 : out <= w[45] ;
	6'b100111 : out <= w[46] ;
	6'b101111 : out <= w[47] ;
	6'b110111 : out <= w[48] ;
	default : out <= 1'bZ;
	endcase
	end
	
endmodule 