
`timescale 1ns/1ns

module tb_lab3_5;


logic out, btn, clk;


detector DUT (.btn(btn), .clk(clk), .out(out));
initial begin
clk = 0;
end
always #1 clk = !clk;
initial begin
btn = 0;
#10 btn = 1;
#1000 btn = 0;
#10 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1000000 btn = 0;
#1000000 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
#1 btn = 0;
#1 btn = 1;
end
initial
#2500000 $stop;

initial begin
$display("Start");

end

endmodule
