module test (p, c);
    
input logic p;
output logic c;

assign c=p

endmodule